�� sr java.util.LinkedList)S]J`�"  xpw   sr model.Memento�'����_� L playert Lmodel/Player;L storaget Lmodel/Storage;xpsr model.PlayerA��6���� I ageI 	eatenFoodI fatnessI 	happinessI hungerI 
meditationI mentalHealthI musclesI physicalHealthI retainedLiquidsI sleepF speedI strengthI trainingChargeI xI yL diseaset Lmodel/Disease;L friendst Ljava/util/ArrayList;L injuryt Lmodel/Injury;L selectedAttacksq ~ L spritest Ljava/util/HashMap;xp   �       P       �    ��������           |                    sr model.Disease�(�l��,� L curesq ~ L effectsq ~ 
L namet Ljava/lang/String;L spriteq ~ L triggersq ~ 
xpsr java.util.ArrayListx����a� I sizexp   w   sr model.actions.MeditationAction&v�p�kp�  xr model.actions.Action�H�ʼE  xpxsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      ~r model.Stats          xr java.lang.Enum          xpt FATNESSsr model.DiseaseInfo�=\E�q�z I pointZ upxp   P~q ~ t MENTAL_HEALTHsq ~   , xt Demenciat demencia.pngsq ~ ?@     w      q ~ sq ~    xsq ~     w    xpsq ~     w    xsq ~ ?@      w       xsr model.Storageu��X@| L 
amountFoodq ~ 
L amountMedicineq ~ 
L foodq ~ 
L medicineq ~ 
xpsq ~ ?@      w       xsq ~ ?@      w       xsq ~ ?@      w       xsq ~ ?@      w       xsq ~ sq ~    �       P       �    ��������           ~                    q ~ q ~ #psq ~     w    xq ~ %sq ~ &q ~ (q ~ )q ~ *q ~ +sq ~ sq ~    �       P       �    ��������           �                    q ~ q ~ #psq ~     w    xq ~ %sq ~ &q ~ (q ~ )q ~ *q ~ +x