�� sr java.util.LinkedList)S]J`�"  xpw   sr model.Memento�'����_� L playert Lmodel/Player;L storaget Lmodel/Storage;xpsr model.PlayerA��6���� I ageI 	eatenFoodI fatnessI 	happinessI hungerI 
meditationI mentalHealthI musclesI physicalHealthI retainedLiquidsI sleepF speedI strengthI trainingChargeI xI yL diseaset Lmodel/Disease;L friendst Ljava/util/ArrayList;L injuryt Lmodel/Injury;L selectedAttacksq ~ L spritest Ljava/util/HashMap;xp      
   P           ������                                sr model.Disease�(�l��,� L curesq ~ L effectsq ~ 
L namet Ljava/lang/String;L spriteq ~ L triggersq ~ 
xpsr java.util.ArrayListx����a� I sizexp   w   sr model.actions.MeditationAction&v�p�kp�  xr model.actions.Action�H�ʼE  xpxsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      ~r model.Stats          xr java.lang.Enum          xpt MENTAL_HEALTHsr model.DiseaseInfo�=\E�q�z I pointZ upxp  , ~q ~ t FATNESSsq ~    Pxt Demenciat demencia.pngsq ~ ?@     w      q ~ sq ~    xsq ~     w    xpsq ~     w    xsq ~ ?@      w       xsr model.Storageu��X@| L 
amountFoodq ~ 
L amountMedicineq ~ 
L foodq ~ 
L medicineq ~ 
xpsq ~ ?@     w      t Galleta Sodasr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp   t Pollo de Pollo landiasq ~ *   t Horpachasq ~ *   t Aguasq ~ *   xsq ~ ?@     w      t Zepolsq ~ *   t Acetaminofensq ~ *   t Paracetamolq ~ 7t TÃ©sq ~ *   
xsq ~ ?@     w      q ~ )sr 
model.Food$g��)I� I energyZ isSolidL nameq ~ xp   q ~ )q ~ -sq ~ <   q ~ -q ~ /sq ~ <   Z q ~ /q ~ 1sq ~ <    q ~ 1xsq ~ ?@     w      q ~ 4sr model.Medicine���!
� I energyL effectsq ~ 
L nameq ~ xp   pq ~ 4q ~ 6sq ~ B   pq ~ 6q ~ 8sq ~ B   sq ~ ?@     w      ~q ~ t STRENGTHsq ~     ~q ~ t HUNGERsq ~    ~q ~ t PHYSICAL_HEALTHsq ~    "q ~ sq ~    xq ~ 8q ~ 9sq ~ B   pq ~ 9xsq ~ sq ~       
   P           ������           &                    q ~ q ~ #psq ~     w    xq ~ %sq ~ &q ~ (q ~ 3q ~ ;q ~ Asq ~ sq ~       
   P           ������           ,                    q ~ q ~ #psq ~     w    xq ~ %sq ~ &q ~ (q ~ 3q ~ ;q ~ Ax