�� sr java.util.LinkedList)S]J`�"  xpw   sr model.Memento�'����_� L playert Lmodel/Player;L storaget Lmodel/Storage;xpsr model.PlayerA��6���� I ageI 	eatenFoodI fatnessI 	happinessI hungerI 
meditationI mentalHealthI musclesI physicalHealthI retainedLiquidsI sleepF speedI strengthI trainingChargeI xI yL diseaset Lmodel/Disease;L friendst Ljava/util/ArrayList;L injuryt Lmodel/Injury;L selectedAttacksq ~ L spritest Ljava/util/HashMap;xp   #      	�       N    ��۬��۬           H                    {sr  java.io.NotSerializableException(Vx �5  xr java.io.ObjectStreamExceptiond��k�9��  xr java.io.IOExceptionl�sde%�  xr java.lang.Exception��>;�  xr java.lang.Throwable��5'9w�� L causet Ljava/lang/Throwable;L detailMessaget Ljava/lang/String;[ 
stackTracet [Ljava/lang/StackTraceElement;L suppressedExceptionst Ljava/util/List;xpq ~ 	t model.Diseaseur [Ljava.lang.StackTraceElement;F*<<�"9  xp   sr java.lang.StackTraceElementa	Ś&6݅ B formatI 
lineNumberL classLoaderNameq ~ L declaringClassq ~ L fileNameq ~ L 
methodNameq ~ L 
moduleNameq ~ L moduleVersionq ~ xp  �pt java.io.ObjectOutputStreamt ObjectOutputStream.javat writeObject0t 	java.baset 11.0.13sq ~   pq ~ q ~ t defaultWriteFieldsq ~ q ~ sq ~   �pq ~ q ~ t writeSerialDataq ~ q ~ sq ~   �pq ~ q ~ t writeOrdinaryObjectq ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   ]pq ~ q ~ t writeObjectq ~ q ~ sq ~   opt java.util.LinkedListt LinkedList.javaq ~  q ~ q ~ sq ~ ����pt -jdk.internal.reflect.GeneratedMethodAccessor6pt invokeq ~ q ~ sq ~    +pt 1jdk.internal.reflect.DelegatingMethodAccessorImplt !DelegatingMethodAccessorImpl.javaq ~ &q ~ q ~ sq ~   6pt java.lang.reflect.Methodt Method.javaq ~ &q ~ q ~ sq ~   ypt java.io.ObjectStreamClasst ObjectStreamClass.javat invokeWriteObjectq ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   ]pq ~ q ~ q ~  q ~ q ~ sq ~    #t appt Utils.MementoReadert MementoReader.javat writeppsq ~    q ~ 6t controller.MementoAdmint MementoAdmin.javat 
addMementoppsq ~    3q ~ 6t controller.ExecutionAdmint ExecutionAdmin.javat runppsq ~   =pt java.lang.Threadt Thread.javaq ~ Aq ~ q ~ sr java.util.Collections$EmptyListz��<���  xpx