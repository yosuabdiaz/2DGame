�� sr java.util.LinkedList)S]J`�"  xpw   sr model.Memento�'����_� L playert Lmodel/Player;L storaget Lmodel/Storage;xpsr model.PlayerA��6���� I ageI 	eatenFoodI fatnessI 	happinessI hungerI 
meditationI mentalHealthI musclesI physicalHealthI retainedLiquidsI sleepF speedI strengthI trainingChargeI xI yL diseaset Lmodel/Disease;L friendst Ljava/util/ArrayList;L injuryt Lmodel/Injury;L selectedAttacksq ~ L spritest Ljava/util/HashMap;xp   2               c                       c                    psr java.util.ArrayListx����a� I sizexp    w    xpsq ~     w    xsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@      w       xsr model.Storage�喩�1� L 
amountFoodq ~ 
L amountMedicineq ~ 
L foodq ~ 
L medicineq ~ 
xpsq ~ ?@      w       xsq ~ ?@      w       xsq ~ ?@      w       xsq ~ ?@      w       xsq ~ sq ~    3               c                       c                    pq ~ psq ~     w    xsq ~ ?@      w       xsq ~ q ~ q ~ q ~ q ~ sq ~ sq ~    4               c                       c                    pq ~ psq ~     w    xsq ~ ?@      w       xsq ~ q ~ q ~ q ~ q ~ sq ~ sq ~    5               c                       c                    pq ~ psq ~     w    xsq ~ ?@      w       xsq ~ q ~ q ~ q ~ q ~ x